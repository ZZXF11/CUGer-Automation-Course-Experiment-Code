library verilog;
use verilog.vl_types.all;
entity xulie_vlg_tst is
end xulie_vlg_tst;
