/*****************文件信息********************************************
**创建日期：   2021.09.08
**版本号：     version 1.0
**功能描述：   按键驱动控制LED
********************************************************************/


module ckey_led(KEY,LEDR);
  input  [3:0] KEY;                   // 四个按键
  output [3:0] LEDR;                  // 四个LED
   
assign LEDR  = KEY;                   //驱动

endmodule